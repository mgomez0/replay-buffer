`timescale 1ns / 1ps
module replay_timer(ack_nack, clk, timer_start);
input ack_nack[1:0];
input clk, timer_start;

